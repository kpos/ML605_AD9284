`timescale 1ns / 1ps

module clock_mgr(
    input clk_in_p,
    input clk_in_n,
    input rst,

    output adc_clk
    );


endmodule
