`timescale 1ns / 1ps

module LVDS_8bit_receiver(input_p[7:0], input_n[7:0], clock_p, clock_n, reset, data[7:0]
    );


endmodule
