`timescale 1ns / 1ps

module test02_top(
    input clk_in_p,
    input clk_in_n,
    input rst,

    input [7:0] adc_data_in_p,
    input [7:0] adc_data_in_n,
    input adc_dco_in_p,
    input adc_dco_in_n,
    output adc_clock_out,
    
    output [7:0] leds,
    output led_C,
    output led_S,
    output led_N
    );

// capture module


 

endmodule


